
module and
(
input a,
input b,
output y
);

y = a & b;
endmodule