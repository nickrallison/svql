module locked_register_async
(
input a,
input b,
output y
);

y = a && b;

endmodule