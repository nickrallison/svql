
module adffe
(
input clk,
input d,
input reset_n,
input en,
output q
);

reg q1;

always @(posedge clk or negedge reset_n) begin
    if (!reset) q1 <= 1'b0;
    else if (en) q1 <= d;
end

assign q = q1;

endmodule